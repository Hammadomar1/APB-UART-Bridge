module DFF(
input x,
input 

  
